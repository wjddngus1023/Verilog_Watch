//MINI_LCD_WATCH.v

module MINI_LCD_WATCH(CLK,RESETN,
LCD_E,LCD_RS,LCD_RW,LCD_DATA,PIEZO,
   KEY1,KEY2,KEY3,KEY4,KEY5,KEY6,KEY7,KEY8);

	input CLK,RESETN;
	input KEY1,KEY2,KEY3,KEY4,KEY5,KEY6,KEY7,KEY8;
	
	output LCD_E, LCD_RS, LCD_RW;
	output [7:0] LCD_DATA;

	wire CLK;
	wire LCD_E, LCD_RS, LCD_RW;
	wire [3:0]H10,H1,M10,M1,S10,S1;

	output PIEZO;
	

	
	
	LCD_WATCH X1(RESETN,CLK,H10,H1,M10,M1,S10,S1,KEY1,KEY2,KEY3,KEY4,KEY5,KEY6,KEY7,KEY8);
	LCD_WATCH_VFD X2(RESETN,CLK,LCD_E, LCD_RS, LCD_RW,LCD_DATA,H10,H1,M10,M1,S10,S1);
	LCD_PIEZO_EX X3(RESETN,CLK,PIEZO);

	
endmodule